module LCD_Controller(reg10_in, segA, segB, segC, segD, segE, segF, segG, an0, dp0);

    input [31:0] reg10_in;
    output wire segA, segB, segC, segD, segE, segF, segG, an0, dp0;

    assign segA = (reg10_in == 32'b00000000000000000000000000000001 || reg10_in == 32'b00000000000000000000000000000100);
    assign segB = (reg10_in == 32'b00000000000000000000000000000101 || reg10_in == 32'b00000000000000000000000000000110);
    assign segC = (reg10_in == 32'b00000000000000000000000000000010);
    assign segD = (reg10_in == 32'b00000000000000000000000000000001 || reg10_in == 32'b00000000000000000000000000000100 || reg10_in == 32'b00000000000000000000000000000111);
    assign segE = (reg10_in == 32'b00000000000000000000000000000001 || reg10_in == 32'b00000000000000000000000000000011 || reg10_in == 32'b00000000000000000000000000000100 || reg10_in == 32'b00000000000000000000000000000101 || reg10_in == 32'b00000000000000000000000000000111 || reg10_in == 32'b00000000000000000000000000001001);
    assign segF = (reg10_in == 32'b00000000000000000000000000000001 || reg10_in == 32'b00000000000000000000000000000010 || reg10_in == 32'b00000000000000000000000000000011 || reg10_in == 32'b00000000000000000000000000000111);
    assign segG = (reg10_in == 32'b00000000000000000000000000000000 || reg10_in == 32'b00000000000000000000000000000001 || reg10_in == 32'b00000000000000000000000000000111);
    assign an0 = 1'b0;
    assign dp0 = 1'b0;


endmodule