module bitwise_not(data_OperandB, result);

    input [31:0] data_OperandB;
    output [31:0] result;

    not result0(result[0], data_OperandB[0]);
    not result1(result[1], data_OperandB[1]);
    not result2(result[2], data_OperandB[2]);
    not result3(result[3], data_OperandB[3]);
    not result4(result[4], data_OperandB[4]);
    not result5(result[5], data_OperandB[5]);
    not result6(result[6], data_OperandB[6]);
    not result7(result[7], data_OperandB[7]);
    not result8(result[8], data_OperandB[8]);
    not result9(result[9], data_OperandB[9]);
    not result10(result[10], data_OperandB[10]);
    not result11(result[11], data_OperandB[11]);
    not result12(result[12], data_OperandB[12]);
    not result13(result[13], data_OperandB[13]);
    not result14(result[14], data_OperandB[14]);
    not result15(result[15], data_OperandB[15]);
    not result16(result[16], data_OperandB[16]);
    not result17(result[17], data_OperandB[17]);
    not result18(result[18], data_OperandB[18]);
    not result19(result[19], data_OperandB[19]);
    not result20(result[20], data_OperandB[20]);
    not result21(result[21], data_OperandB[21]);
    not result22(result[22], data_OperandB[22]);
    not result23(result[23], data_OperandB[23]);
    not result24(result[24], data_OperandB[24]);
    not result25(result[25], data_OperandB[25]);
    not result26(result[26], data_OperandB[26]);
    not result27(result[27], data_OperandB[27]);
    not result28(result[28], data_OperandB[28]);
    not result29(result[29], data_OperandB[29]);
    not result30(result[30], data_OperandB[30]);
    not result31(result[31], data_OperandB[31]);

endmodule